** Profile: "SCHEMATIC1-t"  [ F:\USERS\ROOT\DOCUMENTS\ORCAD\finalvco\t-SCHEMATIC1-t.sim ] 

** Creating circuit file "t-SCHEMATIC1-t.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of F:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1s 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\t-SCHEMATIC1.net" 


.END
